BuzzerRe_inst : BuzzerRe PORT MAP (
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
