library ieee;
use ieee.std_logic_1164.all;

entity map4 is
	port
	(
		F0, F1, F2, F3, F4, F5, F6, F7, F8, F9, F10, F11, F12, F13, F14, F15: out std_logic_vector(31 downto 0)
	);
end map4;	
	
architecture map4_struct of map4 is
begin
	F0 <=  "00100000001000100000110000010000";
	F1 <=  "00000000000000011000110000010000";
	F2 <=  "00010000110000111100000000000000";
	F3 <=  "00000000000000000000001100000000";
	F4 <=  "00010001100100001000001100000000";
	F5 <=  "00000000000000000000001100001000";
	F6 <=  "00010000010000010000000000000000";
	F7 <=  "00000000000000000000000000000010";
	F8 <=  "00000010000010000000110000000000";
	F9 <=  "00000000000001000000110001000100";
	F10 <= "00001100000100110000000000100000";
	F11 <= "00000000001000001000000000000000";
	F12 <= "00000000011000000100000100000010";
	F13 <= "00000010000000000000100000000100";
	F14 <= "00000000010000100000000010000000";
	F15 <= "00010100000010000100010000011000";
end map4_struct;