divisor_inst : divisor PORT MAP (
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
