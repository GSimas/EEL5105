--	ALUNOS:
--	Bruno Luiz da Silva
--	Gustavo Fernades
--
--
--	T�TULO:
--		Expoente
--
--
--	RESUMO:
--		Calcula o expoente baseado na normaliza��o e nos expoentes dados
--
--
--	ENTRADAS/SA�DAS (I/O):
--		(I) a,b: entradas de 4 bits cada que ser�o os expoentes que o usu�rio dar�
--		(I) normal: entrada que receber� o n�mero de vezes que a mantissa foi deslocada para ficar normalizada
--		(I) arguments: argumentos que ser�o recebidos para realizar a soma dos expoentes dados ou o resultado
--					   dessa soma mais o n�mero de deslocamentos realizados.
--		(I) clk,rst: clock e reset, sendo que o reset zera todas sa�das
--		(O) q: sa�da do componente, sendo que ser� esse o expoente final
--
--
--	DESCRI��O:
--		Esse componente ser� respons�vel por dar o expoente da multiplica��o que ser� realizada. Para tal o
--		usu�rio entrar� com os expoentes (em a e b) e dar� o valor "110" para o "argument" para realizar a 
--		soma de ambos. Para previnir casos onde houver uma soma que extrapole o valor "1111" (7 em decimal)
--		ent�o foi adicionado um bit extra na sa�da para armazenar o poss�vel valor extra. Em algum momento
--		ser� enviado o n�mero de deslocamentos realizados para normalizar a mantissa (normal) e assim ter�-se
--		um valor negativo que dever� ser decrementado do atual expoente. Ap�s essa decrementa��o ent�o tem-se
--		o expoente final, por�m ele deve estar na faixa de "0000" a "1111" (0 a 15 em decimal), pois caso
--		extrapole essa faixa ele n�o poder� apresentar o valor correto nos LEDs designados sendo assim um caso
--		de overflow, que ativar� o LED designado para tal.
--
--
--	ANEXO - ARGUMENTS:
--		O "arguments" ser� dado pela FSM e o mesmo � ligado ao bloco de multiplica��o. Aproveitando essa mesma
--		sa�da ent�o usa-se o arguments aqui. Os sinais utilizados e o que fazem s�o:
--
--		110: realiza a soma entre os dois expoentes dados (a e b).
--		111: realiza a subtra��o do atual valor guardado (soma de a e b) com o n�mero de deslocamentos realizados 
--			 na normaliza��o da mantissa.
--
--
--	(I): INPUT	/	(O): OUTPUT

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity expoente is
	generic(N: natural := 4);
	port(
		a,b: in std_logic_vector((N-1) downto 0);		-- Expoentes dados pelo usu�rio
		normal: in std_logic_vector((N-1) downto 0);	-- Deslocamentos que foram necess�rios para normalizar a mantissa
		arguments: in std_logic_vector(2 downto 0);		-- Argumentos que dar� as ordens para o componente
		clk,rst: in std_logic;							-- Clock e reset
		q: out std_logic_vector((N) downto 0)			-- Expoente final
	);
end expoente;

architecture func of expoente is
	signal aux: std_logic_vector(N downto 0);
begin
	EXPOENTE: process(clk,rst)
	begin
		if(rst = '1') then aux <= (others => '0');
		elsif(rising_edge(clk)) then
			if(arguments = "110") then
				-- Soma dos dois expoentes dados com o bit extra para o carry
				aux <= ('0'&a) + ('0'&b);
			elsif(arguments = "111") then
				-- Decremento do resultado da soma anterior com o n�mero de deslocamentos da normaliza��o
				aux <= aux - ('0'&normal);
			else aux <= aux;
			end if;
		end if;
		q <= aux;
	end process;
end func;