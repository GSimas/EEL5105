--	ALUNOS:
--	Bruno Luiz da Silva
--	Gustavo Fernades
--
--
--	T�TULO:
--	Registrador de 16 (+ 1) bits
--
--
--	RESUMO:
--	Registrador de 16 bits com recurso de deslocamento e normaliza��o. � utilizado num multiplicador.
--
--
--	ENTRADAS/SA�DAS (I/O):
--	(I) soma: dado da sa�da do armazenador (soma ou somente a c�pia da parte alta desse registrador)
--	(I) chave: utilizado para carregar a parte baixa do registrador (7 downto 0), sendo conectado nas 
--			   chaves (SW). S� ser� lida quando start tiver valor l�gico alto.
--	(I) start, load: o primeiro ativa a leitura de "chave" e ent�o armazena dados na parte baixa do reg_16.
--					 J� o load permite o armazenamento de "soma" na parte alta do registrador.
--	(I) shift, normalize: recursos extras do registrador que ser�o utilizados para realizar a multiplica��o
--						  de n�meros float. "shift", quando alto, deslocar� os dados para a esquerda
--						  e "normalize" ir� deslocar os dados para a direita e acresentar� 1 ao signal
--						  "exp_aux".
--	(I) clock,reset: clock e reset, sendo que o reset zera todas sa�das
--	(O) q: sa�da dos dados armazenados
-- 	(O) exp: n�mero de vezes em que os dados foram deslocados para direita at� que o LSB fosse 1.
--
--
--	DESCRI��O:
--	Ser�o, primeiramente, dados os valores do multiplicador e estes ser�o guardados na parte baixa do 
--	registrador (7 downto 0). Para tal ser� necess�rio dar um valor l�gico alto para "start".
--	Para carregar o valor que vier do somador ter�-se que colocar um valor l�gico alto em "load" e assim
--	o valor ser� guardado na parte alta do registrador (15 downto 8). 
--
--	Como esse bloco ser� usado para um multiplicador ent�o ser� necess�rio que o valor seja deslocado
--	ap�s a opera��o do componente "somador". Para realizar isto ser� necess�rio dar um valor l�gico alto
--	para "shift" a cada deslocamento desejado.
--
--	A normaliza��o far-se-� necess�ria neste projeto, logo "normalize" deve receber um valor l�gico alto
--	para que inicie-se a normaliza��o. Nesse processo o signal "works" tornar�-se 1 e enquanto o LSB n�o for
--	1, "works" permanecer� em 1, desabilitando qualquer outra opera��o do componente. Quando a opera��o
--	estiver conclu�da ter-se-� o n�mero normalizado e "exp" armazenar� o n�mero de deslocamentos que foram
--	necess�rios.
--
--
--	(I): INPUT	/	(O): OUTPUT

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity reg_16 is 
	port(
		soma: std_logic_vector(8 downto 0);				-- Resultado do somador
		chave: std_logic_vector (7 downto 0);			-- Valor do multiplicador
		start, load, shift, normalize: in std_logic;	-- Recursos para armazenar e manipular valores
		clk, rst: in std_logic;							-- Clock e reset do registrador
		q: out std_logic_vector(15 downto 0);			-- Sa�da (dados armazenados)
		exp: out std_logic_vector(3 downto 0)			-- N�mero de deslocamentos realizados pela normaliza��o
	);
end reg_16;

architecture func of reg_16 is
	signal aux: std_logic_vector(16 downto 0);
	signal exp_aux: std_logic_vector(3 downto 0);
	signal works: std_logic;
begin
	REG16: process(clk,rst)
	begin
		if (rst = '1') then 
			-- Deleta os dados atuais do registrador
			aux <= (others => '0');
			works <= '0';
		elsif (rising_edge(clk)) then 
			if(works = '0') then	
				if(start = '1') then
					-- Carrega o multiplicador para a parte baixa do 
					-- registrador e preenche com 0s a parte alta.
					aux <= '0' & x"00" & chave;
				elsif(load = '1') then
					-- Carrega a soma para a parte baixa do registrador
					aux(16 downto 8) <= soma;
				elsif(shift = '1') then
					-- Desloca os bits uma unidade para a direita.
					aux <= '0' & aux(16 downto 1);
				elsif(normalize = '1') then
					works <= '1';
					exp_aux <= (others => '0');
				end if;
			else 
				if(aux(15) = '0') then
					exp_aux <= exp_aux + 1;
					aux <= aux(15 downto 0) & '0';
				end if;
			end if;
		end if;
		exp <= exp_aux;
		q <= aux(15 downto 0); -- Guarda as opera��es acima efetuadas no registrador.
	end process;
end func;