clock1hz_inst : clock1hz PORT MAP (
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
