divisor5_inst : divisor5 PORT MAP (
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
