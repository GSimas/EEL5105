clockbuzzer1k_inst : clockbuzzer1k PORT MAP (
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
